///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: MUX3
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module testbench();
`include "../Test/Test.v"

///////////////////////////////////////////////////////////////////////////////////
// Inputs: A, B, C (1-bit);  S (2-bit)
reg A, B, C;
reg[1:0] S;
///////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////
// Output: Y (1-bit)
wire Y;
///////////////////////////////////////////////////////////////////////////////////

MUX3 myMUX(.A(A), 
           .B(B), 
           .C(C), 
           .S(S), 
           .Y(Y));

initial begin
////////////////////////////////////////////////////////////////////////////////////////
// Test: S=00
$display("Testing: S=00");
A=1; B=0; C=0; S=2'b00;  #10; 
verifyEqual(Y, A);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: S=01
$display("Testing: S=01");
A=0; B=1; C=0; S=2'b01;  #10; 
verifyEqual(Y, B);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: S=10
$display("Testing: S=10");
A=0; B=0; C=1; S=2'b10;  #10; 
verifyEqual(Y, C);
////////////////////////////////////////////////////////////////////////////////////////

$display("All tests passed.");
end

endmodule